// qsys_core.v

// Generated using ACDS version 15.0 153

`timescale 1 ps / 1 ps
module qsys_core (
		input  wire        avm_cs_i,          //   avm.cs_i
		input  wire [31:0] avm_address_i,     //      .address_i
		input  wire        avm_read_i,        //      .read_i
		output wire        avm_waitrequest_o, //      .waitrequest_o
		output wire [31:0] avm_readdata_o,    //      .readdata_o
		input  wire        avm_write_i,       //      .write_i
		input  wire [31:0] avm_writedata_i,   //      .writedata_i
		input  wire [3:0]  avm_byteenable_i,  //      .byteenable_i
		input  wire        clk_clk,           //   clk.clk
		input  wire        reset_reset_n,     // reset.reset_n
		output wire [12:0] sdram_addr,        // sdram.addr
		output wire [1:0]  sdram_ba,          //      .ba
		output wire        sdram_cas_n,       //      .cas_n
		output wire        sdram_cke,         //      .cke
		output wire        sdram_cs_n,        //      .cs_n
		inout  wire [15:0] sdram_dq,          //      .dq
		output wire [1:0]  sdram_dqm,         //      .dqm
		output wire        sdram_ras_n,       //      .ras_n
		output wire        sdram_we_n         //      .we_n
	);

	wire         wb_avm_bridge_m0_chipselect;              // wb_avm_bridge:avm_cs -> mm_interconnect_0:wb_avm_bridge_m0_chipselect
	wire         wb_avm_bridge_m0_waitrequest;             // mm_interconnect_0:wb_avm_bridge_m0_waitrequest -> wb_avm_bridge:avm_waitrequest
	wire  [31:0] wb_avm_bridge_m0_readdata;                // mm_interconnect_0:wb_avm_bridge_m0_readdata -> wb_avm_bridge:avm_readdata
	wire  [31:0] wb_avm_bridge_m0_address;                 // wb_avm_bridge:avm_address -> mm_interconnect_0:wb_avm_bridge_m0_address
	wire         wb_avm_bridge_m0_read;                    // wb_avm_bridge:avm_read -> mm_interconnect_0:wb_avm_bridge_m0_read
	wire   [3:0] wb_avm_bridge_m0_byteenable;              // wb_avm_bridge:avm_byteenable -> mm_interconnect_0:wb_avm_bridge_m0_byteenable
	wire         wb_avm_bridge_m0_write;                   // wb_avm_bridge:avm_write -> mm_interconnect_0:wb_avm_bridge_m0_write
	wire  [31:0] wb_avm_bridge_m0_writedata;               // wb_avm_bridge:avm_writedata -> mm_interconnect_0:wb_avm_bridge_m0_writedata
	wire         mm_interconnect_0_sdram_s1_chipselect;    // mm_interconnect_0:sdram_s1_chipselect -> sdram:az_cs
	wire  [15:0] mm_interconnect_0_sdram_s1_readdata;      // sdram:za_data -> mm_interconnect_0:sdram_s1_readdata
	wire         mm_interconnect_0_sdram_s1_waitrequest;   // sdram:za_waitrequest -> mm_interconnect_0:sdram_s1_waitrequest
	wire  [24:0] mm_interconnect_0_sdram_s1_address;       // mm_interconnect_0:sdram_s1_address -> sdram:az_addr
	wire         mm_interconnect_0_sdram_s1_read;          // mm_interconnect_0:sdram_s1_read -> sdram:az_rd_n
	wire   [1:0] mm_interconnect_0_sdram_s1_byteenable;    // mm_interconnect_0:sdram_s1_byteenable -> sdram:az_be_n
	wire         mm_interconnect_0_sdram_s1_readdatavalid; // sdram:za_valid -> mm_interconnect_0:sdram_s1_readdatavalid
	wire         mm_interconnect_0_sdram_s1_write;         // mm_interconnect_0:sdram_s1_write -> sdram:az_wr_n
	wire  [15:0] mm_interconnect_0_sdram_s1_writedata;     // mm_interconnect_0:sdram_s1_writedata -> sdram:az_data

	qsys_core_sdram sdram (
		.clk            (clk_clk),                                  //   clk.clk
		.reset_n        (reset_reset_n),                            // reset.reset_n
		.az_addr        (mm_interconnect_0_sdram_s1_address),       //    s1.address
		.az_be_n        (~mm_interconnect_0_sdram_s1_byteenable),   //      .byteenable_n
		.az_cs          (mm_interconnect_0_sdram_s1_chipselect),    //      .chipselect
		.az_data        (mm_interconnect_0_sdram_s1_writedata),     //      .writedata
		.az_rd_n        (~mm_interconnect_0_sdram_s1_read),         //      .read_n
		.az_wr_n        (~mm_interconnect_0_sdram_s1_write),        //      .write_n
		.za_data        (mm_interconnect_0_sdram_s1_readdata),      //      .readdata
		.za_valid       (mm_interconnect_0_sdram_s1_readdatavalid), //      .readdatavalid
		.za_waitrequest (mm_interconnect_0_sdram_s1_waitrequest),   //      .waitrequest
		.zs_addr        (sdram_addr),                               //  wire.export
		.zs_ba          (sdram_ba),                                 //      .export
		.zs_cas_n       (sdram_cas_n),                              //      .export
		.zs_cke         (sdram_cke),                                //      .export
		.zs_cs_n        (sdram_cs_n),                               //      .export
		.zs_dq          (sdram_dq),                                 //      .export
		.zs_dqm         (sdram_dqm),                                //      .export
		.zs_ras_n       (sdram_ras_n),                              //      .export
		.zs_we_n        (sdram_we_n)                                //      .export
	);

	wb_avm_bridge_if wb_avm_bridge (
		.clk             (clk_clk),                      //   clock.clk
		.reset           (~reset_reset_n),               //   reset.reset
		.avm_cs          (wb_avm_bridge_m0_chipselect),  //      m0.chipselect
		.avm_address     (wb_avm_bridge_m0_address),     //        .address
		.avm_read        (wb_avm_bridge_m0_read),        //        .read
		.avm_waitrequest (wb_avm_bridge_m0_waitrequest), //        .waitrequest
		.avm_readdata    (wb_avm_bridge_m0_readdata),    //        .readdata
		.avm_write       (wb_avm_bridge_m0_write),       //        .write
		.avm_writedata   (wb_avm_bridge_m0_writedata),   //        .writedata
		.avm_byteenable  (wb_avm_bridge_m0_byteenable),  //        .byteenable
		.cs_i            (avm_cs_i),                     // conduit.cs_i
		.address_i       (avm_address_i),                //        .address_i
		.read_i          (avm_read_i),                   //        .read_i
		.waitrequest_o   (avm_waitrequest_o),            //        .waitrequest_o
		.readdata_o      (avm_readdata_o),               //        .readdata_o
		.write_i         (avm_write_i),                  //        .write_i
		.writedata_i     (avm_writedata_i),              //        .writedata_i
		.byteenable_i    (avm_byteenable_i)              //        .byteenable_i
	);

	qsys_core_mm_interconnect_0 mm_interconnect_0 (
		.clk_sys_clk_clk                                 (clk_clk),                                  //                               clk_sys_clk.clk
		.wb_avm_bridge_reset_reset_bridge_in_reset_reset (~reset_reset_n),                           // wb_avm_bridge_reset_reset_bridge_in_reset.reset
		.wb_avm_bridge_m0_address                        (wb_avm_bridge_m0_address),                 //                          wb_avm_bridge_m0.address
		.wb_avm_bridge_m0_waitrequest                    (wb_avm_bridge_m0_waitrequest),             //                                          .waitrequest
		.wb_avm_bridge_m0_byteenable                     (wb_avm_bridge_m0_byteenable),              //                                          .byteenable
		.wb_avm_bridge_m0_chipselect                     (wb_avm_bridge_m0_chipselect),              //                                          .chipselect
		.wb_avm_bridge_m0_read                           (wb_avm_bridge_m0_read),                    //                                          .read
		.wb_avm_bridge_m0_readdata                       (wb_avm_bridge_m0_readdata),                //                                          .readdata
		.wb_avm_bridge_m0_write                          (wb_avm_bridge_m0_write),                   //                                          .write
		.wb_avm_bridge_m0_writedata                      (wb_avm_bridge_m0_writedata),               //                                          .writedata
		.sdram_s1_address                                (mm_interconnect_0_sdram_s1_address),       //                                  sdram_s1.address
		.sdram_s1_write                                  (mm_interconnect_0_sdram_s1_write),         //                                          .write
		.sdram_s1_read                                   (mm_interconnect_0_sdram_s1_read),          //                                          .read
		.sdram_s1_readdata                               (mm_interconnect_0_sdram_s1_readdata),      //                                          .readdata
		.sdram_s1_writedata                              (mm_interconnect_0_sdram_s1_writedata),     //                                          .writedata
		.sdram_s1_byteenable                             (mm_interconnect_0_sdram_s1_byteenable),    //                                          .byteenable
		.sdram_s1_readdatavalid                          (mm_interconnect_0_sdram_s1_readdatavalid), //                                          .readdatavalid
		.sdram_s1_waitrequest                            (mm_interconnect_0_sdram_s1_waitrequest),   //                                          .waitrequest
		.sdram_s1_chipselect                             (mm_interconnect_0_sdram_s1_chipselect)     //                                          .chipselect
	);

endmodule
